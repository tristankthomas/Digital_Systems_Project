`define CLK_PERIOD_ns   20